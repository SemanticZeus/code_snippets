* 


E1 1 0 2 3 5
R1 1 2 1
R2 1 3 10
I1 0 2 10
R3 2 3 2
G1 3 0 1 3 .1

.tran 1m 1

.control
run
plot v(1)-v(2) v(1) v(2) v(3)
.endc
.end

