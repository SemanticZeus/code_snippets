* VCO
.model npn npn(BF=300)

.MODEL BC547BP NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5
+IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80
+VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33

.include "modelos_subckt/ti/ua741.mod"

vin vin 0 sin (5 5 1)
VDC vcc 0 10
VDC2 0 vee 5
R1 vin vn 100k
R2 vin vp 50k
C1 vn output_opamp1 .1u ic=0

* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |

X1 vp vn vcc vee output_opamp1 UA741 
Rshort1 output_opamp1 triangle_output 0
Rshort2 output_opamp1 vn2 0
R4 vn 2 50k
VIC1 2 tr1c 0
R3 vp 0 50k

* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |

X2 vp2 vn2 vcc vee output_opamp2 UA741
R6 vp2 output_opamp2 100k
Rshort3 output_opamp2 square_output 0
R7 vp2 0 100k
R8 vcc vp2 100k
R5 output_opamp2 tr1b 220



Q1 tr1c tr1b 0 npn

.tran 10u 2 uic

.control
run
plot v(square_output) v(triangle_output) 

.endc
.end
