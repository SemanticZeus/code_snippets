



V1 1 0 1
R1 1 0 1k


G1 0 2  1 0 2
RL 2 0 1

.tran 1m 1

.control
run
plot v(1) v(2)
.endc
.end

