* simulating key in ngspice

.MODEL BC546 NPN (IS=50.7F NF=1 BF=318 VAF=145 IKF=.3
+ ISE=15.9P NE=2 BR=4 NR=1 VAR=24 IKR=.45 RE=1.54 RB=6.17
+ RC=.617 XTB=1.5 CJE=20.8P CJC=8.33P TF=611P TR=138N)
*   National 65 Volt  .5 Amp  260 MHz  SiNPN  Transistor  01-26-1991
*PINOUT TO-92 3 2 1


.SUBCKT KEY in node1 node2
Q1 collectoro base emitter BC546
RE emitter GND


