*FM foster seeley Discriminator Circuit



V1 in 0 SFFM(0 10 100k 5 10.7MEG)
Rs in 1 0
C1 1 0 13.3p
L1 1 0 17.6u
L2 2 m1 8.8u
L3 m1 3 8.8u
K1 L1 L2 .222
K2 L1 L3 .222

Cc 1 m1 10u

C2 2 3 13.3pf
R3 2 3 10k
D1 2 a1 diode
D2 3 a2 diode
R1 a1 m2 1000
R2 a2 m2 1000
C3 a1 m2 .1u
C4 a2 m2 .1u
Lrfc m1 m2 1u
CL a1 a2 .1u
RL a1 a2 10k
Rshort1 a2 0 0
*Rshort2 m2 0 0

.tran 1n 10m

.model diode D(Is=1e-10 n=1e-3)

.control
run
plot v(a1)

.endc

.end
