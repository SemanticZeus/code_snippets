* ideal diode

.MODEL DI_1N4001G D  ( IS=65.4p RS=4.2m BV=5000.0 IBV=5.00u
+ CJO=14.8p  M=0.333 N=1.36 TT=2.88u )

.subckt ideal_diode anode cathod

E1 out1 0 vp1 vn1 100
D1 out1 o1 DI_1N4001G

Rshort1 anode vp1 0
RShort2 o1 vn1 0

Rshort3 o1 cathod 0

.ends


V1 1 0 sin(0 1 1)
X1 1 2 ideal_diode
R1 2 0 1k

D1 1 3 DI_1N4001G
R2 3 0 1k

 
.tran 100u 5 uic

.control
run
plot V(1) V(2) V(3)
.endc
.end
