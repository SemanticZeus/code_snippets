* Ideal Diode Example Circuit

V1 Vin 0 sin(0 5 10)        ; 5V DC source
R1 Vin Anode 1k      ; Series resistor
D1 Anode Cathode D_ideal
RL Cathode 0 1k      ; Load resistor

.model D_ideal D (IS=1e-15 N=0.01 RS=1e-6 TT=0 CJO=0 EG=1e6 BV=1e9 IBV=1e-3)

.control
  tran 1m 1        ; Transient analysis from 0 to 10µs
  plot V(Anode) V(Cathode) v(Vin)
.endc
.end
